`include "multibank_memory.sv"